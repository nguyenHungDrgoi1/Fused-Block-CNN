module top_module (
    input clk,
    input rst_n,
    
);
endmodule