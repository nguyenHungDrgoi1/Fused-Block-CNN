module PE_4mul (
    input wire          clk,
    input wire          en,

    input wire [7:0]    IFM1, IFM2, IFM3, IFM4,
    input wire [7:0]    Weight1, Weight2, Weight3, Weight4,

    
);
endmodule